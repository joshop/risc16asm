typedef enum logic [3:0] { NAND, AND, NOR, OR, ADD, SUB, XOR, SL, SR } alu_func_e;
