typedef logic [3:0] enum {
  NAND,
  AND,
  NOR,
  OR,
  ADD,
  SUB,
  XOR,
  SL,
  SR
} alu_func_e;
