typedef enum logic [2:0] { OPIMM, OP, LUI, BRANCH, JALR, LOAD, STORE } itype_e;
// typedef enum logic [3:0] { NAND, AND, NOR, OR, ADD, SUB, XOR, SL, SR } alu_func_e;
// typedef enum logic [2:0] { BZ, BNZ, BP, BNP } br_func_e;
